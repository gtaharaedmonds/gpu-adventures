module rgb2dvi (
    output logic tsms
);


endmodule
